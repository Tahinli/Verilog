module hello_world;
    initial begin
        $display ("Hello World");
        $finish;
    end
endmodule